 1  ||   Vitello tonnato    ;   15    ||       Antipasto misto ;   15    ||      Riso col nero di seppie ;    16        ||      Ossobuco  ; 25      ||   Panna cotta ;   7     ||     Aqua  ; 10   ||       Te nero   ;   4     ||      Spuma  ;  4    
   2  ||   Vitello tonnato  ;  15,67   ||   Orechiette pugliesi con salsiccia toscana piccante    ;  17     ||      Panna cotta  ;  7     ||     Caffe freddo    ;    5    ||   Spuma  ; 4   ||       Aqua  ; 10  


  3   ||    Insalata mista  ;   8,99       ||    Antipasto misto   ;    15        ||       Saltimboca   ;   17        ||   Cappon magro  ;  28   ||    Panna cotta   ;    7        ||     Te nero ; 4    

 4   ||   Vitello tonnato ;   15      ||     Insalata frutti di mare    ; 15     ||     Saltimboca   ;  17     ||   Tirami su  ;    8  ||    Cappucino   ;  4        ||    Espresso   ;   4  ||   Cappucino  ;    4    

 5   ||    Insalata Caprese ;  10      ||   Arrosto di manzo   ;  25   ||   Tirami su  ; 8       ||    Aqua ; 10    ||    Spuma ;  4    


   6  ||  Antipasto misto  ; 15        ||     Insalata mista    ; 8   ||   Saltimboca ;    17     ||  Pizza Margerita    ;  12   ||     Marsala-Zabaione ;   6    ||     Marsala-Zabaione  ;    6    ||    Espresso  ;   4     ||    Coca  ;  3     ||     Cappucino  ; 4 


 7  ||   Insalata mista   ;  8      ||      Insalata mista   ;  8   ||     Penne arrabiata    ;    15      ||     Caffe freddo ; 5        ||      Cappucino  ;  4     ||       Cappucino ;   4  



   8 ||    Antipasto misto  ;  15       ||       Cozze al marinara  ;   16       ||      Tirami su    ;  8      ||    Panna cotta  ;   7    ||      Aqua  ;   10   

    9 ||  Vitello tonnato  ;    15       ||       Ossobuco    ;  25   ||     Marsala-Zabaione   ;    6      ||   Espresso    ; 4  


    10    ||   Insalata Caprese    ;  10        ||      Saltimboca  ;    17  ||    Scallopine al limone   ;  27     ||      Caffe freddo  ; 5  ||      Espresso   ;  4   ||   Espresso   ;    4    ||        Aqua  ;   10   

